-------------------------------------------------------------------------------------------
--    ▄▄   ▄▄ ▄▄▄▄▄▄ ▄▄▄     ▄▄▄▄▄▄▄    ▄▄▄▄▄▄▄ ▄▄▄▄▄▄  ▄▄▄▄▄▄  ▄▄▄▄▄▄▄ ▄▄▄▄▄▄   
--   █  █ █  █      █   █   █       █  █       █      ██      ██       █   ▄  █  
--   █  █▄█  █  ▄   █   █   █    ▄▄▄█  █   ▄   █  ▄    █  ▄    █    ▄▄▄█  █ █ █  
--   █       █ █▄█  █   █   █   █▄▄▄   █  █▄█  █ █ █   █ █ █   █   █▄▄▄█   █▄▄█▄ 
--   █   ▄   █      █   █▄▄▄█    ▄▄▄█  █       █ █▄█   █ █▄█   █    ▄▄▄█    ▄▄  █
--   █  █ █  █  ▄   █       █   █      █   ▄   █       █       █   █▄▄▄█   █  █ █
--   █▄▄█ █▄▄█▄█ █▄▄█▄▄▄▄▄▄▄█▄▄▄█      █▄▄█ █▄▄█▄▄▄▄▄▄██▄▄▄▄▄▄██▄▄▄▄▄▄▄█▄▄▄█  █▄█
-- ________________________________________________________________________________________
-- @author. LathiasMaar
-- @brief. This code implements a half_adder circuit
-- 
-- @components. Xor2 gates, And2 gates, Or2 gates
--
-- @function. if (a xor b) = 1:         
--                sum = 1;                        
--            else:                                        
--                sum = 0;                            
--                                                          
--            if (a and b):                    
--                car = 1;                        
--            else :                      
--                car = 0;
--
-- @truth_table.
--      _______________________
--    /|  A  |  B  | Out | CAR |
--   | | --- | --- | --- | --- |          Inputs                Outputs
--   | |  0  |  0  |  0  |  0  |                   ___________
--   | |  1  |  0  |  1  |  0  |                  |           \
--   | |  0  |  1  |  1  |  0  |             A ---|  H_ADDER  |-- Sum 
--   | |  1  |  1  |  0  |  1  |             B ---|___________|-- Car  
--   |/ ¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯/
--    ¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯¯
-------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;

library libs;
use libs.all;
-------------------------------------------------------------------------------------------
entity HalfAdder is
    PORT(
        a, b : IN std_logic;
        sum, car : OUT std_logic
    );
end HalfAdder;
-------------------------------------------------------------------------------------------
architecture structure of HalfAdder is

    component Xor2 is
        PORT(
            a,b : IN std_logic;
            y : OUT std_logic
        );   
    end component;

    component And2
        PORT(
            a,b : IN std_logic;
            y : OUT std_logic);
    end component;

    begin
        U1: Xor2 PORT map(
            a => a,
            b => b,
            y => sum     
        );

        U2: And2 PORT map(
            a => a,
            b => b,
            y => car  
        );
end structure;
-------------------------------------------------------------------------------------------